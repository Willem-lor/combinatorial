// Code your design here
module mux2 ();

endmodule


module mux4 ();

endmodule


module mux8 ();

endmodule


module adder ();

endmodule


module multiplier ();

endmodule


module alu ();

endmodule
